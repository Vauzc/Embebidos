`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:42:43 05/04/2020 
// Design Name: 
// Module Name:    osf 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module osf(
    input in,
    output M1L,
    output M1R,
    output M1O,
    output M2L,
    output M2R,
    output M2O,
    output M3L,
    output M3R,
    output M3O,
    output M4L,
    output M4R,
    output M4O
    );


endmodule
